`timescale 1ns/1ps
module ROM(addr,data);
input [30:0] addr;
output reg [31:0] data;
wire [28:0] index;
assign index=addr[30:2];
always @(*)
begin
  case(index)
  0:data<=32'b00001000000000000000000000000011;
  1:data<=32'b00001000000000000000000000110101;
  2:data<=32'b00001000000000000000000010000100;
  3:data<=32'b00110000000111010000000000000000;
  4:data<=32'b00111100000100000100000000000000;
  5:data<=32'b00000000000000001000100000100111;
  6:data<=32'b10101110000000000000000000001000;
  7:data<=32'b10101110000000000000000000001100;
  8:data<=32'b00100000000010000000011111111111;
  9:data<=32'b10101110000010000000000000010100;
  10:data<=32'b00100000000010000000000000000011;
  11:data<=32'b10101110000010000000000000100000;
  12:data<=32'b10101110000100010000000000000100;
  13:data<=32'b00100010001010001000101011010000;
  14:data<=32'b00100001000010001000101011010000;
  15:data<=32'b10101110000010000000000000000000;
  16:data<=32'b00100000000010000000000000000011;
  17:data<=32'b10101110000010000000000000001000;
  18:data<=32'b00100000000100100000000000000010;
  19:data<=32'b10001110000010000000000000100000;
  20:data<=32'b00110001000010010000000000001100;
  21:data<=32'b00000000000010010100100011000010;
  22:data<=32'b00011001001000001111111111111100;
  23:data<=32'b00100010010100101111111111111111;
  24:data<=32'b00011010010000000000000000000010;
  25:data<=32'b10001110000001000000000000011100;
  26:data<=32'b00001000000000000000000000010011;
  27:data<=32'b00100000000100100000000000000010;
  28:data<=32'b10001110000001010000000000011100;
  29:data<=32'b00000000100000000011000000100000;
  30:data<=32'b00000000101000000011100000100000;
  31:data<=32'b00000000110001110100100000101010;
  32:data<=32'b00010101001000000000000000000011;
  33:data<=32'b00000000000001100100000000100000;
  34:data<=32'b00000000000001110011000000100000;
  35:data<=32'b00000000000010000011100000100000;
  36:data<=32'b00000000111001100011100000100010;
  37:data<=32'b00000000110001110100100000101010;
  38:data<=32'b00010101001000001111111111111101;
  39:data<=32'b00010000111000000000000000000101;
  40:data<=32'b00000000000000000000000000000000;
  41:data<=32'b00000000000001100100000000100000;
  42:data<=32'b00000000000001110011000000100000;
  43:data<=32'b00000000000010000011100000100000;
  44:data<=32'b00001000000000000000000000100100;
  45:data<=32'b00000000000001100001000000100000;
  46:data<=32'b10101110000000100000000000001100;
  47:data<=32'b10001110000010000000000000100000;
  48:data<=32'b00110001000010010000000000010000;
  49:data<=32'b00000000000010010100100100000010;
  50:data<=32'b00010101001000001111111111111100;
  51:data<=32'b10101110000000100000000000011000;
  52:data<=32'b00001000000000000000000000010011;
  53:data<=32'b10001110000110010000000000001000;
  54:data<=32'b00110011001110010000000000000001;
  55:data<=32'b10101110000110010000000000001000;
  56:data<=32'b00000001000000001001100000100000;
  57:data<=32'b00000001001000001010000000100000;
  58:data<=32'b10001110000010000000000000010100;
  59:data<=32'b00110001000010010000111100000000;
  60:data<=32'b00100000000010100000011100000000;
  61:data<=32'b00010101001010100000000000000011;
  62:data<=32'b00100000000010010000101100000000;
  63:data<=32'b00110000100010110000000000001111;
  64:data<=32'b00001000000000000000000001001111;
  65:data<=32'b00100000000010100000101100000000;
  66:data<=32'b00010101001010100000000000000100;
  67:data<=32'b00100000000010010000110100000000;
  68:data<=32'b00110000101010110000000011110000;
  69:data<=32'b00000000000010110101100100000010;
  70:data<=32'b00001000000000000000000001001111;
  71:data<=32'b00100000000010100000110100000000;
  72:data<=32'b00010101001010100000000000000011;
  73:data<=32'b00100000000010010000111000000000;
  74:data<=32'b00110000101010110000000000001111;
  75:data<=32'b00001000000000000000000001001111;
  76:data<=32'b00100000000010010000011100000000;
  77:data<=32'b00110000100010110000000011110000;
  78:data<=32'b00000000000010110101100100000010;
  79:data<=32'b00100000000011000000000011000000;
  80:data<=32'b00011001011000000000000000101011;
  81:data<=32'b00100001011010111111111111111111;
  82:data<=32'b00100000000011000000000011111001;
  83:data<=32'b00011001011000000000000000101000;
  84:data<=32'b00100001011010111111111111111111;
  85:data<=32'b00100000000011000000000010100100;
  86:data<=32'b00011001011000000000000000100101;
  87:data<=32'b00100001011010111111111111111111;
  88:data<=32'b00100000000011000000000010110000;
  89:data<=32'b00011001011000000000000000100010;
  90:data<=32'b00100001011010111111111111111111;
  91:data<=32'b00100000000011000000000010011001;
  92:data<=32'b00011001011000000000000000011111;
  93:data<=32'b00100001011010111111111111111111;
  94:data<=32'b00100000000011000000000010010010;
  95:data<=32'b00011001011000000000000000011100;
  96:data<=32'b00100001011010111111111111111111;
  97:data<=32'b00100000000011000000000010000010;
  98:data<=32'b00011001011000000000000000011001;
  99:data<=32'b00100001011010111111111111111111;
  100:data<=32'b00100000000011000000000011111000;
  101:data<=32'b00011001011000000000000000010110;
  102:data<=32'b00100001011010111111111111111111;
  103:data<=32'b00100000000011000000000010000000;
  104:data<=32'b00011001011000000000000000010011;
  105:data<=32'b00100001011010111111111111111111;
  106:data<=32'b00100000000011000000000010010000;
  107:data<=32'b00011001011000000000000000010000;
  108:data<=32'b00100001011010111111111111111111;
  109:data<=32'b00100000000011000000000010001000;
  110:data<=32'b00011001011000000000000000001101;
  111:data<=32'b00100001011010111111111111111111;
  112:data<=32'b00100000000011000000000010000011;
  113:data<=32'b00011001011000000000000000001010;
  114:data<=32'b00100001011010111111111111111111;
  115:data<=32'b00100000000011000000000011000110;
  116:data<=32'b00011001011000000000000000000111;
  117:data<=32'b00100001011010111111111111111111;
  118:data<=32'b00100000000011000000000010100001;
  119:data<=32'b00011001011000000000000000000100;
  120:data<=32'b00100001011010111111111111111111;
  121:data<=32'b00100000000011000000000010000110;
  122:data<=32'b00011001011000000000000000000001;
  123:data<=32'b00100000000011000000000010001110;
  124:data<=32'b00000001001011000100000000100101;
  125:data<=32'b10101110000010000000000000010100;
  126:data<=32'b00000010011000000100000000100000;
  127:data<=32'b00000010100000000100100000100000;
  128:data<=32'b10001110000110010000000000001000;
  129:data<=32'b00110111001110010000000000000010;
  130:data<=32'b10101110000110010000000000001000;
  131:data<=32'b00000011010000000000000000001000;
  132:data<=32'b00100000000010000000011100000000;
  133:data<=32'b10101110000010000000000000010100;
  134:data<=32'b00001000000000000000000010000100;
default:data<=32'hffffffff;
endcase

end

endmodule



